`ifndef _ct_vh_
`define _ct_vh_

`define RESET_VAL 1
`timescale 1ns / 1ps

`endif
`ifndef _ct_vh_
`define _ct_vh_

`define RESET_VAL 1
`define INT_SIZE 8

`define WIDTH_IN 8
`define WIDTH_OUT 8
`define N_LLRS 4
`define EXTENDED_BITS 4
`define N_V 31
`define E 140
`define N_ITER 5
`define CROSS_P 0.01

`timescale 1ns / 1ps

`endif
`timescale 1ns / 1ps
`define RESET_VAL 1

module variable_nodes
	#(  parameter WIDTH = 8,
	    parameter N_V = 31,
	    parameter E = 140)
	( input clk, rst,
	  input data_ready,
	  input prev_ready,
	  input [WIDTH * N_V - 1 : 0] all_llrs,
	  input [WIDTH * E - 1 : 0] prev_proc_elem,
	  output [WIDTH * E - 1 : 0] proc_elem,
	  output reg varn_ready);

	localparam EXTENDED_WIDTH = WIDTH + 4;
	reg [EXTENDED_WIDTH * E - 1 : 0] temp_reg, temp_reg_nxt;

	saturate #(.WIDTH(WIDTH), .EXTENDED_BITS(EXTENDED_WIDTH - WIDTH)) sat[E - 1 : 0] (.in(temp_reg), .out(proc_elem));

	always @(posedge clk) begin
		if (rst == `RESET_VAL) begin
			varn_ready <= 1'b0;
		end
		else if (prev_ready == 1 && data_ready == 1) begin
			temp_reg <= temp_reg_nxt;

			varn_ready <= 1'b1;
		end
	end

	always @* begin
		temp_reg_nxt = temp_reg;

		if (prev_ready == 1 && data_ready == 1) begin
			temp_reg_nxt[(EXTENDED_WIDTH * 1) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 1) - 1]}}, all_llrs[(WIDTH * 1) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 1) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 1) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 2) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 1) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 1) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 3) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 1) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 1) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 4) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 1) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 1) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 5) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 1) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 1) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 6) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 1) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 1) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 7) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 1) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 1) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 8) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 1) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 1) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 9) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 1) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 1) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 10) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 2) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 1) - 1]}}, all_llrs[(WIDTH * 1) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 2) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 2) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 1) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 2) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 2) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 3) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 2) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 2) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 4) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 2) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 2) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 5) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 2) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 2) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 6) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 2) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 2) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 7) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 2) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 2) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 8) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 2) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 2) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 9) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 2) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 2) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 10) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 3) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 1) - 1]}}, all_llrs[(WIDTH * 1) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 3) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 3) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 1) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 3) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 3) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 2) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 3) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 3) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 4) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 3) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 3) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 5) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 3) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 3) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 6) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 3) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 3) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 7) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 3) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 3) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 8) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 3) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 3) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 9) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 3) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 3) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 10) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 4) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 1) - 1]}}, all_llrs[(WIDTH * 1) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 4) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 4) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 1) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 4) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 4) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 2) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 4) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 4) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 3) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 4) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 4) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 5) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 4) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 4) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 6) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 4) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 4) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 7) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 4) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 4) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 8) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 4) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 4) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 9) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 4) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 4) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 10) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 5) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 1) - 1]}}, all_llrs[(WIDTH * 1) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 5) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 5) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 1) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 5) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 5) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 2) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 5) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 5) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 3) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 5) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 5) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 4) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 5) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 5) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 6) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 5) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 5) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 7) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 5) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 5) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 8) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 5) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 5) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 9) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 5) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 5) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 10) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 6) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 1) - 1]}}, all_llrs[(WIDTH * 1) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 6) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 6) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 1) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 6) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 6) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 2) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 6) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 6) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 3) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 6) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 6) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 4) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 6) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 6) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 5) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 6) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 6) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 7) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 6) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 6) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 8) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 6) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 6) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 9) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 6) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 6) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 10) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 7) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 1) - 1]}}, all_llrs[(WIDTH * 1) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 7) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 7) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 1) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 7) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 7) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 2) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 7) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 7) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 3) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 7) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 7) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 4) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 7) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 7) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 5) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 7) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 7) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 6) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 7) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 7) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 8) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 7) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 7) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 9) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 7) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 7) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 10) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 8) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 1) - 1]}}, all_llrs[(WIDTH * 1) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 8) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 8) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 1) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 8) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 8) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 2) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 8) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 8) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 3) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 8) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 8) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 4) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 8) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 8) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 5) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 8) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 8) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 6) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 8) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 8) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 7) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 8) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 8) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 9) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 8) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 8) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 10) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 9) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 1) - 1]}}, all_llrs[(WIDTH * 1) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 9) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 9) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 1) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 9) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 9) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 2) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 9) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 9) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 3) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 9) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 9) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 4) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 9) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 9) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 5) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 9) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 9) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 6) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 9) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 9) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 7) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 9) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 9) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 8) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 9) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 9) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 10) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 10) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 1) - 1]}}, all_llrs[(WIDTH * 1) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 10) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 10) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 1) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 10) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 10) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 2) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 10) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 10) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 3) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 10) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 10) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 4) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 10) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 10) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 5) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 10) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 10) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 6) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 10) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 10) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 7) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 10) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 10) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 8) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 10) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 10) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 9) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 11) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 2) - 1]}}, all_llrs[(WIDTH * 2) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 11) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 11) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 12) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 11) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 11) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 13) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 11) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 11) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 14) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 11) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 11) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 15) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 11) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 11) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 16) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 11) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 11) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 17) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 12) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 2) - 1]}}, all_llrs[(WIDTH * 2) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 12) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 12) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 11) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 12) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 12) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 13) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 12) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 12) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 14) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 12) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 12) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 15) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 12) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 12) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 16) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 12) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 12) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 17) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 13) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 2) - 1]}}, all_llrs[(WIDTH * 2) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 13) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 13) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 11) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 13) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 13) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 12) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 13) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 13) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 14) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 13) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 13) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 15) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 13) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 13) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 16) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 13) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 13) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 17) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 14) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 2) - 1]}}, all_llrs[(WIDTH * 2) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 14) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 14) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 11) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 14) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 14) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 12) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 14) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 14) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 13) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 14) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 14) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 15) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 14) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 14) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 16) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 14) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 14) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 17) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 15) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 2) - 1]}}, all_llrs[(WIDTH * 2) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 15) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 15) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 11) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 15) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 15) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 12) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 15) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 15) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 13) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 15) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 15) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 14) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 15) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 15) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 16) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 15) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 15) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 17) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 16) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 2) - 1]}}, all_llrs[(WIDTH * 2) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 16) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 16) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 11) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 16) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 16) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 12) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 16) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 16) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 13) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 16) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 16) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 14) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 16) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 16) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 15) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 16) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 16) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 17) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 17) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 2) - 1]}}, all_llrs[(WIDTH * 2) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 17) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 17) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 11) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 17) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 17) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 12) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 17) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 17) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 13) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 17) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 17) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 14) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 17) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 17) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 15) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 17) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 17) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 16) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 18) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 3) - 1]}}, all_llrs[(WIDTH * 3) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 18) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 18) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 19) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 18) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 18) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 20) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 18) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 18) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 21) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 18) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 18) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 22) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 18) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 18) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 23) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 18) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 18) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 24) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 19) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 3) - 1]}}, all_llrs[(WIDTH * 3) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 19) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 19) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 18) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 19) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 19) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 20) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 19) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 19) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 21) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 19) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 19) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 22) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 19) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 19) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 23) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 19) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 19) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 24) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 20) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 3) - 1]}}, all_llrs[(WIDTH * 3) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 20) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 20) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 18) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 20) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 20) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 19) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 20) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 20) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 21) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 20) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 20) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 22) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 20) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 20) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 23) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 20) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 20) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 24) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 21) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 3) - 1]}}, all_llrs[(WIDTH * 3) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 21) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 21) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 18) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 21) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 21) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 19) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 21) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 21) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 20) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 21) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 21) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 22) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 21) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 21) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 23) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 21) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 21) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 24) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 22) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 3) - 1]}}, all_llrs[(WIDTH * 3) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 22) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 22) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 18) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 22) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 22) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 19) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 22) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 22) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 20) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 22) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 22) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 21) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 22) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 22) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 23) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 22) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 22) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 24) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 23) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 3) - 1]}}, all_llrs[(WIDTH * 3) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 23) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 23) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 18) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 23) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 23) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 19) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 23) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 23) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 20) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 23) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 23) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 21) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 23) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 23) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 22) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 23) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 23) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 24) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 24) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 3) - 1]}}, all_llrs[(WIDTH * 3) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 24) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 24) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 18) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 24) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 24) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 19) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 24) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 24) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 20) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 24) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 24) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 21) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 24) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 24) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 22) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 24) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 24) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 23) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 25) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 4) - 1]}}, all_llrs[(WIDTH * 4) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 25) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 25) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 26) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 25) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 25) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 27) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 25) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 25) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 28) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 25) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 25) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 29) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 25) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 25) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 30) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 25) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 25) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 31) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 26) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 4) - 1]}}, all_llrs[(WIDTH * 4) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 26) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 26) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 25) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 26) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 26) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 27) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 26) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 26) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 28) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 26) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 26) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 29) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 26) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 26) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 30) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 26) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 26) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 31) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 27) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 4) - 1]}}, all_llrs[(WIDTH * 4) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 27) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 27) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 25) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 27) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 27) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 26) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 27) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 27) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 28) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 27) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 27) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 29) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 27) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 27) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 30) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 27) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 27) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 31) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 28) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 4) - 1]}}, all_llrs[(WIDTH * 4) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 28) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 28) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 25) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 28) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 28) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 26) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 28) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 28) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 27) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 28) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 28) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 29) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 28) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 28) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 30) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 28) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 28) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 31) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 29) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 4) - 1]}}, all_llrs[(WIDTH * 4) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 29) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 29) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 25) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 29) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 29) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 26) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 29) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 29) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 27) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 29) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 29) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 28) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 29) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 29) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 30) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 29) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 29) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 31) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 30) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 4) - 1]}}, all_llrs[(WIDTH * 4) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 30) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 30) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 25) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 30) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 30) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 26) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 30) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 30) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 27) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 30) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 30) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 28) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 30) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 30) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 29) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 30) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 30) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 31) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 31) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 4) - 1]}}, all_llrs[(WIDTH * 4) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 31) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 31) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 25) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 31) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 31) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 26) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 31) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 31) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 27) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 31) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 31) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 28) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 31) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 31) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 29) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 31) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 31) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 30) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 32) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 5) - 1]}}, all_llrs[(WIDTH * 5) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 32) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 32) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 33) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 32) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 32) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 34) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 32) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 32) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 35) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 32) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 32) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 36) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 32) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 32) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 37) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 33) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 5) - 1]}}, all_llrs[(WIDTH * 5) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 33) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 33) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 32) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 33) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 33) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 34) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 33) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 33) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 35) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 33) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 33) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 36) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 33) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 33) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 37) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 34) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 5) - 1]}}, all_llrs[(WIDTH * 5) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 34) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 34) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 32) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 34) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 34) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 33) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 34) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 34) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 35) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 34) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 34) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 36) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 34) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 34) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 37) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 35) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 5) - 1]}}, all_llrs[(WIDTH * 5) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 35) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 35) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 32) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 35) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 35) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 33) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 35) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 35) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 34) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 35) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 35) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 36) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 35) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 35) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 37) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 36) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 5) - 1]}}, all_llrs[(WIDTH * 5) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 36) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 36) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 32) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 36) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 36) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 33) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 36) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 36) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 34) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 36) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 36) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 35) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 36) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 36) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 37) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 37) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 5) - 1]}}, all_llrs[(WIDTH * 5) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 37) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 37) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 32) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 37) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 37) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 33) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 37) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 37) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 34) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 37) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 37) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 35) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 37) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 37) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 36) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 38) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 6) - 1]}}, all_llrs[(WIDTH * 6) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 38) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 38) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 39) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 38) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 38) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 40) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 38) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 38) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 41) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 38) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 38) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 42) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 38) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 38) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 43) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 39) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 6) - 1]}}, all_llrs[(WIDTH * 6) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 39) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 39) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 38) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 39) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 39) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 40) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 39) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 39) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 41) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 39) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 39) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 42) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 39) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 39) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 43) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 40) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 6) - 1]}}, all_llrs[(WIDTH * 6) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 40) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 40) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 38) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 40) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 40) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 39) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 40) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 40) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 41) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 40) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 40) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 42) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 40) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 40) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 43) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 41) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 6) - 1]}}, all_llrs[(WIDTH * 6) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 41) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 41) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 38) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 41) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 41) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 39) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 41) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 41) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 40) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 41) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 41) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 42) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 41) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 41) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 43) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 42) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 6) - 1]}}, all_llrs[(WIDTH * 6) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 42) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 42) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 38) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 42) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 42) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 39) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 42) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 42) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 40) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 42) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 42) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 41) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 42) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 42) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 43) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 43) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 6) - 1]}}, all_llrs[(WIDTH * 6) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 43) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 43) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 38) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 43) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 43) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 39) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 43) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 43) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 40) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 43) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 43) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 41) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 43) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 43) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 42) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 44) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 7) - 1]}}, all_llrs[(WIDTH * 7) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 44) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 44) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 45) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 44) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 44) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 46) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 44) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 44) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 47) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 44) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 44) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 48) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 44) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 44) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 49) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 45) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 7) - 1]}}, all_llrs[(WIDTH * 7) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 45) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 45) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 44) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 45) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 45) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 46) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 45) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 45) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 47) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 45) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 45) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 48) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 45) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 45) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 49) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 46) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 7) - 1]}}, all_llrs[(WIDTH * 7) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 46) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 46) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 44) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 46) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 46) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 45) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 46) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 46) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 47) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 46) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 46) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 48) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 46) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 46) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 49) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 47) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 7) - 1]}}, all_llrs[(WIDTH * 7) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 47) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 47) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 44) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 47) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 47) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 45) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 47) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 47) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 46) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 47) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 47) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 48) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 47) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 47) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 49) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 48) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 7) - 1]}}, all_llrs[(WIDTH * 7) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 48) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 48) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 44) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 48) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 48) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 45) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 48) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 48) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 46) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 48) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 48) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 47) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 48) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 48) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 49) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 49) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 7) - 1]}}, all_llrs[(WIDTH * 7) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 49) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 49) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 44) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 49) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 49) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 45) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 49) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 49) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 46) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 49) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 49) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 47) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 49) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 49) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 48) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 50) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 8) - 1]}}, all_llrs[(WIDTH * 8) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 50) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 50) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 51) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 50) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 50) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 52) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 50) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 50) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 53) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 50) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 50) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 54) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 50) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 50) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 55) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 51) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 8) - 1]}}, all_llrs[(WIDTH * 8) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 51) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 51) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 50) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 51) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 51) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 52) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 51) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 51) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 53) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 51) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 51) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 54) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 51) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 51) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 55) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 52) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 8) - 1]}}, all_llrs[(WIDTH * 8) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 52) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 52) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 50) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 52) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 52) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 51) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 52) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 52) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 53) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 52) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 52) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 54) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 52) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 52) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 55) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 53) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 8) - 1]}}, all_llrs[(WIDTH * 8) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 53) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 53) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 50) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 53) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 53) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 51) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 53) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 53) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 52) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 53) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 53) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 54) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 53) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 53) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 55) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 54) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 8) - 1]}}, all_llrs[(WIDTH * 8) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 54) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 54) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 50) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 54) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 54) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 51) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 54) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 54) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 52) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 54) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 54) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 53) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 54) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 54) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 55) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 55) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 8) - 1]}}, all_llrs[(WIDTH * 8) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 55) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 55) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 50) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 55) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 55) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 51) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 55) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 55) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 52) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 55) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 55) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 53) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 55) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 55) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 54) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 56) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 9) - 1]}}, all_llrs[(WIDTH * 9) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 56) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 56) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 57) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 56) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 56) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 58) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 56) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 56) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 59) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 56) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 56) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 60) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 56) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 56) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 61) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 57) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 9) - 1]}}, all_llrs[(WIDTH * 9) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 57) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 57) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 56) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 57) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 57) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 58) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 57) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 57) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 59) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 57) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 57) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 60) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 57) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 57) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 61) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 58) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 9) - 1]}}, all_llrs[(WIDTH * 9) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 58) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 58) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 56) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 58) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 58) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 57) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 58) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 58) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 59) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 58) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 58) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 60) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 58) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 58) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 61) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 59) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 9) - 1]}}, all_llrs[(WIDTH * 9) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 59) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 59) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 56) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 59) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 59) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 57) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 59) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 59) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 58) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 59) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 59) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 60) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 59) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 59) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 61) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 60) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 9) - 1]}}, all_llrs[(WIDTH * 9) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 60) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 60) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 56) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 60) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 60) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 57) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 60) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 60) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 58) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 60) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 60) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 59) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 60) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 60) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 61) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 61) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 9) - 1]}}, all_llrs[(WIDTH * 9) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 61) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 61) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 56) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 61) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 61) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 57) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 61) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 61) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 58) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 61) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 61) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 59) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 61) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 61) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 60) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 62) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 10) - 1]}}, all_llrs[(WIDTH * 10) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 62) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 62) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 63) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 62) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 62) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 64) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 62) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 62) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 65) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 62) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 62) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 66) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 62) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 62) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 67) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 62) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 62) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 68) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 63) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 10) - 1]}}, all_llrs[(WIDTH * 10) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 63) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 63) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 62) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 63) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 63) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 64) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 63) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 63) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 65) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 63) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 63) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 66) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 63) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 63) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 67) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 63) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 63) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 68) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 64) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 10) - 1]}}, all_llrs[(WIDTH * 10) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 64) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 64) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 62) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 64) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 64) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 63) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 64) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 64) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 65) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 64) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 64) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 66) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 64) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 64) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 67) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 64) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 64) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 68) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 65) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 10) - 1]}}, all_llrs[(WIDTH * 10) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 65) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 65) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 62) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 65) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 65) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 63) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 65) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 65) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 64) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 65) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 65) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 66) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 65) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 65) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 67) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 65) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 65) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 68) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 66) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 10) - 1]}}, all_llrs[(WIDTH * 10) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 66) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 66) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 62) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 66) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 66) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 63) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 66) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 66) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 64) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 66) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 66) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 65) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 66) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 66) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 67) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 66) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 66) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 68) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 67) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 10) - 1]}}, all_llrs[(WIDTH * 10) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 67) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 67) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 62) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 67) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 67) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 63) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 67) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 67) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 64) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 67) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 67) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 65) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 67) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 67) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 66) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 67) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 67) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 68) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 68) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 10) - 1]}}, all_llrs[(WIDTH * 10) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 68) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 68) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 62) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 68) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 68) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 63) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 68) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 68) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 64) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 68) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 68) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 65) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 68) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 68) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 66) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 68) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 68) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 67) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 69) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 11) - 1]}}, all_llrs[(WIDTH * 11) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 69) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 69) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 70) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 69) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 69) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 71) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 69) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 69) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 72) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 69) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 69) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 73) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 69) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 69) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 74) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 70) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 11) - 1]}}, all_llrs[(WIDTH * 11) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 70) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 70) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 69) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 70) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 70) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 71) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 70) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 70) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 72) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 70) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 70) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 73) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 70) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 70) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 74) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 71) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 11) - 1]}}, all_llrs[(WIDTH * 11) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 71) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 71) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 69) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 71) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 71) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 70) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 71) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 71) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 72) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 71) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 71) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 73) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 71) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 71) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 74) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 72) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 11) - 1]}}, all_llrs[(WIDTH * 11) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 72) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 72) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 69) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 72) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 72) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 70) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 72) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 72) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 71) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 72) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 72) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 73) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 72) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 72) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 74) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 73) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 11) - 1]}}, all_llrs[(WIDTH * 11) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 73) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 73) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 69) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 73) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 73) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 70) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 73) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 73) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 71) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 73) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 73) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 72) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 73) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 73) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 74) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 74) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 11) - 1]}}, all_llrs[(WIDTH * 11) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 74) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 74) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 69) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 74) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 74) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 70) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 74) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 74) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 71) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 74) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 74) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 72) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 74) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 74) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 73) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 75) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 12) - 1]}}, all_llrs[(WIDTH * 12) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 75) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 75) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 76) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 75) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 75) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 77) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 75) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 75) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 78) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 75) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 75) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 79) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 75) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 75) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 80) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 75) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 75) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 81) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 75) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 75) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 82) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 75) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 75) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 83) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 75) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 75) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 84) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 75) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 75) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 85) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 76) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 12) - 1]}}, all_llrs[(WIDTH * 12) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 76) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 76) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 75) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 76) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 76) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 77) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 76) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 76) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 78) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 76) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 76) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 79) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 76) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 76) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 80) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 76) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 76) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 81) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 76) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 76) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 82) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 76) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 76) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 83) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 76) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 76) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 84) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 76) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 76) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 85) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 77) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 12) - 1]}}, all_llrs[(WIDTH * 12) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 77) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 77) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 75) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 77) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 77) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 76) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 77) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 77) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 78) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 77) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 77) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 79) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 77) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 77) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 80) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 77) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 77) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 81) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 77) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 77) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 82) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 77) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 77) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 83) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 77) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 77) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 84) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 77) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 77) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 85) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 78) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 12) - 1]}}, all_llrs[(WIDTH * 12) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 78) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 78) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 75) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 78) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 78) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 76) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 78) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 78) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 77) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 78) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 78) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 79) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 78) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 78) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 80) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 78) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 78) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 81) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 78) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 78) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 82) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 78) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 78) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 83) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 78) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 78) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 84) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 78) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 78) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 85) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 79) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 12) - 1]}}, all_llrs[(WIDTH * 12) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 79) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 79) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 75) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 79) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 79) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 76) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 79) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 79) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 77) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 79) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 79) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 78) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 79) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 79) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 80) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 79) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 79) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 81) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 79) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 79) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 82) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 79) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 79) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 83) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 79) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 79) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 84) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 79) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 79) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 85) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 80) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 12) - 1]}}, all_llrs[(WIDTH * 12) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 80) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 80) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 75) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 80) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 80) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 76) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 80) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 80) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 77) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 80) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 80) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 78) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 80) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 80) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 79) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 80) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 80) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 81) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 80) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 80) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 82) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 80) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 80) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 83) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 80) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 80) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 84) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 80) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 80) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 85) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 81) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 12) - 1]}}, all_llrs[(WIDTH * 12) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 81) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 81) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 75) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 81) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 81) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 76) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 81) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 81) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 77) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 81) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 81) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 78) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 81) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 81) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 79) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 81) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 81) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 80) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 81) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 81) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 82) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 81) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 81) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 83) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 81) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 81) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 84) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 81) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 81) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 85) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 82) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 12) - 1]}}, all_llrs[(WIDTH * 12) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 82) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 82) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 75) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 82) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 82) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 76) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 82) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 82) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 77) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 82) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 82) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 78) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 82) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 82) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 79) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 82) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 82) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 80) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 82) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 82) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 81) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 82) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 82) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 83) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 82) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 82) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 84) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 82) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 82) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 85) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 83) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 12) - 1]}}, all_llrs[(WIDTH * 12) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 83) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 83) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 75) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 83) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 83) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 76) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 83) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 83) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 77) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 83) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 83) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 78) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 83) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 83) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 79) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 83) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 83) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 80) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 83) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 83) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 81) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 83) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 83) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 82) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 83) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 83) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 84) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 83) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 83) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 85) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 84) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 12) - 1]}}, all_llrs[(WIDTH * 12) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 84) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 84) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 75) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 84) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 84) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 76) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 84) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 84) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 77) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 84) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 84) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 78) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 84) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 84) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 79) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 84) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 84) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 80) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 84) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 84) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 81) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 84) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 84) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 82) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 84) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 84) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 83) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 84) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 84) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 85) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 85) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 12) - 1]}}, all_llrs[(WIDTH * 12) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 85) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 85) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 75) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 85) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 85) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 76) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 85) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 85) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 77) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 85) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 85) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 78) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 85) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 85) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 79) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 85) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 85) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 80) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 85) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 85) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 81) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 85) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 85) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 82) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 85) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 85) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 83) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 85) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 85) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 84) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 86) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 13) - 1]}}, all_llrs[(WIDTH * 13) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 86) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 86) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 87) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 86) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 86) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 88) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 86) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 86) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 89) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 86) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 86) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 90) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 86) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 86) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 91) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 86) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 86) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 92) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 86) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 86) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 93) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 86) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 86) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 94) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 86) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 86) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 95) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 87) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 13) - 1]}}, all_llrs[(WIDTH * 13) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 87) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 87) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 86) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 87) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 87) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 88) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 87) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 87) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 89) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 87) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 87) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 90) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 87) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 87) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 91) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 87) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 87) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 92) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 87) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 87) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 93) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 87) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 87) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 94) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 87) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 87) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 95) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 88) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 13) - 1]}}, all_llrs[(WIDTH * 13) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 88) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 88) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 86) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 88) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 88) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 87) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 88) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 88) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 89) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 88) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 88) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 90) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 88) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 88) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 91) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 88) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 88) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 92) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 88) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 88) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 93) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 88) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 88) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 94) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 88) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 88) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 95) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 89) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 13) - 1]}}, all_llrs[(WIDTH * 13) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 89) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 89) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 86) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 89) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 89) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 87) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 89) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 89) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 88) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 89) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 89) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 90) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 89) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 89) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 91) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 89) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 89) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 92) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 89) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 89) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 93) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 89) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 89) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 94) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 89) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 89) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 95) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 90) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 13) - 1]}}, all_llrs[(WIDTH * 13) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 90) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 90) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 86) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 90) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 90) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 87) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 90) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 90) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 88) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 90) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 90) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 89) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 90) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 90) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 91) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 90) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 90) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 92) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 90) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 90) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 93) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 90) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 90) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 94) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 90) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 90) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 95) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 91) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 13) - 1]}}, all_llrs[(WIDTH * 13) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 91) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 91) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 86) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 91) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 91) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 87) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 91) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 91) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 88) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 91) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 91) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 89) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 91) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 91) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 90) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 91) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 91) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 92) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 91) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 91) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 93) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 91) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 91) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 94) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 91) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 91) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 95) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 92) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 13) - 1]}}, all_llrs[(WIDTH * 13) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 92) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 92) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 86) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 92) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 92) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 87) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 92) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 92) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 88) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 92) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 92) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 89) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 92) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 92) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 90) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 92) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 92) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 91) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 92) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 92) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 93) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 92) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 92) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 94) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 92) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 92) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 95) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 93) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 13) - 1]}}, all_llrs[(WIDTH * 13) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 93) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 93) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 86) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 93) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 93) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 87) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 93) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 93) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 88) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 93) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 93) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 89) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 93) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 93) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 90) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 93) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 93) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 91) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 93) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 93) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 92) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 93) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 93) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 94) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 93) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 93) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 95) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 94) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 13) - 1]}}, all_llrs[(WIDTH * 13) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 94) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 94) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 86) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 94) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 94) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 87) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 94) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 94) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 88) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 94) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 94) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 89) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 94) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 94) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 90) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 94) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 94) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 91) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 94) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 94) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 92) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 94) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 94) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 93) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 94) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 94) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 95) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 95) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 13) - 1]}}, all_llrs[(WIDTH * 13) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 95) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 95) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 86) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 95) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 95) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 87) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 95) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 95) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 88) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 95) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 95) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 89) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 95) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 95) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 90) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 95) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 95) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 91) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 95) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 95) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 92) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 95) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 95) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 93) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 95) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 95) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 94) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 96) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 14) - 1]}}, all_llrs[(WIDTH * 14) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 96) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 96) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 97) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 96) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 96) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 98) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 96) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 96) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 99) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 96) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 96) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 100) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 96) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 96) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 101) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 96) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 96) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 102) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 96) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 96) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 103) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 96) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 96) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 104) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 96) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 96) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 105) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 97) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 14) - 1]}}, all_llrs[(WIDTH * 14) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 97) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 97) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 96) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 97) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 97) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 98) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 97) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 97) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 99) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 97) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 97) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 100) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 97) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 97) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 101) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 97) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 97) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 102) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 97) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 97) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 103) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 97) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 97) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 104) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 97) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 97) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 105) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 98) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 14) - 1]}}, all_llrs[(WIDTH * 14) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 98) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 98) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 96) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 98) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 98) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 97) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 98) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 98) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 99) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 98) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 98) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 100) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 98) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 98) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 101) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 98) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 98) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 102) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 98) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 98) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 103) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 98) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 98) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 104) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 98) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 98) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 105) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 99) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 14) - 1]}}, all_llrs[(WIDTH * 14) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 99) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 99) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 96) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 99) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 99) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 97) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 99) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 99) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 98) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 99) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 99) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 100) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 99) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 99) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 101) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 99) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 99) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 102) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 99) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 99) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 103) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 99) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 99) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 104) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 99) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 99) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 105) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 100) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 14) - 1]}}, all_llrs[(WIDTH * 14) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 100) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 100) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 96) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 100) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 100) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 97) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 100) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 100) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 98) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 100) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 100) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 99) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 100) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 100) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 101) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 100) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 100) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 102) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 100) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 100) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 103) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 100) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 100) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 104) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 100) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 100) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 105) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 101) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 14) - 1]}}, all_llrs[(WIDTH * 14) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 101) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 101) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 96) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 101) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 101) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 97) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 101) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 101) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 98) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 101) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 101) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 99) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 101) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 101) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 100) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 101) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 101) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 102) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 101) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 101) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 103) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 101) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 101) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 104) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 101) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 101) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 105) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 102) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 14) - 1]}}, all_llrs[(WIDTH * 14) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 102) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 102) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 96) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 102) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 102) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 97) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 102) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 102) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 98) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 102) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 102) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 99) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 102) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 102) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 100) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 102) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 102) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 101) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 102) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 102) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 103) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 102) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 102) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 104) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 102) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 102) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 105) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 103) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 14) - 1]}}, all_llrs[(WIDTH * 14) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 103) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 103) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 96) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 103) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 103) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 97) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 103) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 103) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 98) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 103) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 103) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 99) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 103) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 103) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 100) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 103) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 103) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 101) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 103) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 103) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 102) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 103) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 103) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 104) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 103) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 103) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 105) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 104) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 14) - 1]}}, all_llrs[(WIDTH * 14) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 104) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 104) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 96) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 104) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 104) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 97) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 104) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 104) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 98) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 104) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 104) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 99) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 104) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 104) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 100) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 104) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 104) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 101) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 104) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 104) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 102) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 104) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 104) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 103) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 104) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 104) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 105) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 105) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 14) - 1]}}, all_llrs[(WIDTH * 14) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 105) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 105) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 96) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 105) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 105) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 97) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 105) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 105) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 98) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 105) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 105) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 99) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 105) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 105) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 100) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 105) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 105) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 101) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 105) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 105) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 102) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 105) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 105) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 103) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 105) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 105) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 104) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 106) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 15) - 1]}}, all_llrs[(WIDTH * 15) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 106) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 106) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 107) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 106) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 106) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 108) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 106) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 106) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 109) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 106) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 106) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 110) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 106) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 106) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 111) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 106) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 106) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 112) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 106) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 106) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 113) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 106) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 106) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 114) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 106) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 106) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 115) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 107) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 15) - 1]}}, all_llrs[(WIDTH * 15) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 107) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 107) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 106) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 107) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 107) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 108) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 107) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 107) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 109) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 107) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 107) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 110) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 107) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 107) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 111) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 107) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 107) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 112) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 107) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 107) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 113) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 107) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 107) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 114) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 107) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 107) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 115) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 108) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 15) - 1]}}, all_llrs[(WIDTH * 15) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 108) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 108) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 106) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 108) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 108) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 107) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 108) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 108) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 109) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 108) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 108) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 110) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 108) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 108) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 111) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 108) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 108) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 112) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 108) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 108) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 113) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 108) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 108) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 114) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 108) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 108) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 115) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 109) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 15) - 1]}}, all_llrs[(WIDTH * 15) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 109) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 109) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 106) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 109) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 109) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 107) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 109) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 109) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 108) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 109) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 109) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 110) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 109) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 109) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 111) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 109) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 109) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 112) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 109) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 109) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 113) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 109) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 109) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 114) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 109) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 109) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 115) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 110) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 15) - 1]}}, all_llrs[(WIDTH * 15) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 110) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 110) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 106) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 110) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 110) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 107) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 110) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 110) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 108) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 110) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 110) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 109) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 110) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 110) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 111) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 110) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 110) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 112) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 110) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 110) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 113) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 110) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 110) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 114) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 110) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 110) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 115) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 111) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 15) - 1]}}, all_llrs[(WIDTH * 15) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 111) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 111) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 106) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 111) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 111) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 107) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 111) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 111) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 108) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 111) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 111) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 109) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 111) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 111) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 110) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 111) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 111) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 112) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 111) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 111) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 113) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 111) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 111) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 114) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 111) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 111) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 115) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 112) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 15) - 1]}}, all_llrs[(WIDTH * 15) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 112) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 112) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 106) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 112) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 112) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 107) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 112) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 112) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 108) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 112) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 112) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 109) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 112) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 112) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 110) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 112) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 112) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 111) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 112) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 112) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 113) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 112) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 112) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 114) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 112) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 112) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 115) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 113) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 15) - 1]}}, all_llrs[(WIDTH * 15) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 113) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 113) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 106) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 113) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 113) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 107) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 113) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 113) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 108) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 113) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 113) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 109) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 113) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 113) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 110) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 113) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 113) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 111) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 113) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 113) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 112) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 113) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 113) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 114) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 113) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 113) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 115) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 114) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 15) - 1]}}, all_llrs[(WIDTH * 15) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 114) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 114) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 106) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 114) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 114) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 107) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 114) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 114) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 108) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 114) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 114) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 109) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 114) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 114) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 110) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 114) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 114) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 111) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 114) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 114) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 112) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 114) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 114) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 113) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 114) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 114) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 115) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 115) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 15) - 1]}}, all_llrs[(WIDTH * 15) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 115) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 115) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 106) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 115) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 115) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 107) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 115) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 115) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 108) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 115) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 115) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 109) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 115) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 115) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 110) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 115) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 115) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 111) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 115) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 115) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 112) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 115) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 115) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 113) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 115) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 115) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 114) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 116) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 16) - 1]}}, all_llrs[(WIDTH * 16) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 116) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 116) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 117) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 116) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 116) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 118) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 116) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 116) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 119) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 116) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 116) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 120) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 116) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 116) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 121) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 116) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 116) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 122) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 116) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 116) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 123) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 116) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 116) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 124) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 116) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 116) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 125) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 117) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 16) - 1]}}, all_llrs[(WIDTH * 16) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 117) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 117) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 116) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 117) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 117) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 118) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 117) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 117) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 119) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 117) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 117) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 120) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 117) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 117) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 121) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 117) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 117) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 122) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 117) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 117) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 123) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 117) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 117) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 124) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 117) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 117) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 125) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 118) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 16) - 1]}}, all_llrs[(WIDTH * 16) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 118) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 118) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 116) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 118) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 118) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 117) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 118) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 118) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 119) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 118) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 118) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 120) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 118) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 118) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 121) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 118) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 118) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 122) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 118) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 118) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 123) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 118) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 118) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 124) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 118) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 118) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 125) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 119) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 16) - 1]}}, all_llrs[(WIDTH * 16) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 119) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 119) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 116) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 119) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 119) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 117) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 119) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 119) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 118) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 119) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 119) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 120) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 119) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 119) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 121) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 119) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 119) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 122) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 119) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 119) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 123) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 119) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 119) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 124) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 119) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 119) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 125) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 120) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 16) - 1]}}, all_llrs[(WIDTH * 16) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 120) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 120) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 116) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 120) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 120) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 117) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 120) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 120) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 118) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 120) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 120) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 119) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 120) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 120) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 121) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 120) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 120) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 122) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 120) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 120) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 123) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 120) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 120) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 124) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 120) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 120) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 125) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 121) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 16) - 1]}}, all_llrs[(WIDTH * 16) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 121) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 121) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 116) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 121) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 121) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 117) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 121) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 121) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 118) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 121) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 121) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 119) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 121) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 121) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 120) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 121) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 121) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 122) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 121) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 121) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 123) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 121) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 121) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 124) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 121) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 121) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 125) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 122) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 16) - 1]}}, all_llrs[(WIDTH * 16) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 122) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 122) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 116) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 122) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 122) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 117) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 122) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 122) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 118) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 122) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 122) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 119) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 122) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 122) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 120) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 122) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 122) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 121) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 122) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 122) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 123) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 122) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 122) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 124) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 122) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 122) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 125) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 123) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 16) - 1]}}, all_llrs[(WIDTH * 16) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 123) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 123) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 116) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 123) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 123) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 117) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 123) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 123) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 118) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 123) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 123) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 119) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 123) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 123) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 120) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 123) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 123) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 121) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 123) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 123) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 122) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 123) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 123) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 124) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 123) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 123) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 125) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 124) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 16) - 1]}}, all_llrs[(WIDTH * 16) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 124) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 124) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 116) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 124) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 124) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 117) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 124) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 124) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 118) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 124) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 124) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 119) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 124) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 124) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 120) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 124) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 124) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 121) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 124) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 124) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 122) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 124) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 124) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 123) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 124) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 124) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 125) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 125) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 16) - 1]}}, all_llrs[(WIDTH * 16) - 1 -: WIDTH]};
			temp_reg_nxt[(EXTENDED_WIDTH * 125) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 125) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 116) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 125) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 125) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 117) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 125) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 125) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 118) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 125) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 125) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 119) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 125) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 125) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 120) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 125) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 125) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 121) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 125) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 125) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 122) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 125) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 125) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 123) - 1 -: WIDTH];
			temp_reg_nxt[(EXTENDED_WIDTH * 125) - 1 -: EXTENDED_WIDTH] = temp_reg_nxt[(EXTENDED_WIDTH * 125) - 1 -: EXTENDED_WIDTH] + prev_proc_elem[(WIDTH * 124) - 1 -: WIDTH];

			temp_reg_nxt[(EXTENDED_WIDTH * 126) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 17) - 1]}}, all_llrs[(WIDTH * 17) - 1 -: WIDTH]};

			temp_reg_nxt[(EXTENDED_WIDTH * 127) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 18) - 1]}}, all_llrs[(WIDTH * 18) - 1 -: WIDTH]};

			temp_reg_nxt[(EXTENDED_WIDTH * 128) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 19) - 1]}}, all_llrs[(WIDTH * 19) - 1 -: WIDTH]};

			temp_reg_nxt[(EXTENDED_WIDTH * 129) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 20) - 1]}}, all_llrs[(WIDTH * 20) - 1 -: WIDTH]};

			temp_reg_nxt[(EXTENDED_WIDTH * 130) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 21) - 1]}}, all_llrs[(WIDTH * 21) - 1 -: WIDTH]};

			temp_reg_nxt[(EXTENDED_WIDTH * 131) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 22) - 1]}}, all_llrs[(WIDTH * 22) - 1 -: WIDTH]};

			temp_reg_nxt[(EXTENDED_WIDTH * 132) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 23) - 1]}}, all_llrs[(WIDTH * 23) - 1 -: WIDTH]};

			temp_reg_nxt[(EXTENDED_WIDTH * 133) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 24) - 1]}}, all_llrs[(WIDTH * 24) - 1 -: WIDTH]};

			temp_reg_nxt[(EXTENDED_WIDTH * 134) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 25) - 1]}}, all_llrs[(WIDTH * 25) - 1 -: WIDTH]};

			temp_reg_nxt[(EXTENDED_WIDTH * 135) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 26) - 1]}}, all_llrs[(WIDTH * 26) - 1 -: WIDTH]};

			temp_reg_nxt[(EXTENDED_WIDTH * 136) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 27) - 1]}}, all_llrs[(WIDTH * 27) - 1 -: WIDTH]};

			temp_reg_nxt[(EXTENDED_WIDTH * 137) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 28) - 1]}}, all_llrs[(WIDTH * 28) - 1 -: WIDTH]};

			temp_reg_nxt[(EXTENDED_WIDTH * 138) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 29) - 1]}}, all_llrs[(WIDTH * 29) - 1 -: WIDTH]};

			temp_reg_nxt[(EXTENDED_WIDTH * 139) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 30) - 1]}}, all_llrs[(WIDTH * 30) - 1 -: WIDTH]};

			temp_reg_nxt[(EXTENDED_WIDTH * 140) - 1 -: EXTENDED_WIDTH] = {{(EXTENDED_WIDTH - WIDTH){all_llrs[(WIDTH * 31) - 1]}}, all_llrs[(WIDTH * 31) - 1 -: WIDTH]};

		end
	end
endmodule
